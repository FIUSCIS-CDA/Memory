///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: RAM (CLK=200)
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020, 2025 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module testbenchRAM();
`include "../Test/Test.v"

//////////////////////////////////////////////////////////////////////////////////
// Tests both synchronous and asynchronous memory
/////////////////////////////////////////////////////////////
// Inputs: addr, writedata (32-bit), we (1-bit)
//         clk (1-bit, synchronous only)
reg[31:0] addr;
reg[31:0] writedata;
reg we;
reg clk; // Clock it at 200
/////////////////////////////////////////////////////////////
// Outputs: readdataSynch (32-bit, synchronous only)
wire[31:0] readdataSynch;
/////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////

RAM DMemorySynch(
	.clk(clk),
	.a(addr),
	.rd(readdataSynch),
        .wd(writedata),
        .we(we));


initial begin
/////////////////////////////////////////////////////////////////////////////
// Populate both memories with the same data
$readmemh("datamem.dat",DMemorySynch.memory);
/////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////
// For both memories, address 8 has the value 2 initially
////////////////////////////////////////////////////////////////////////////
// Test: addr=8, writedata=42, we=0 (readdata should still be 2)
addr=8; we=0; writedata=42; #100;
$display("[SYNCH] Testing addr=8 with writedata=42 and we=0: DM[8]=2"); 
verifyEqual32(readdataSynch, 2);
///////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////
// Test: addr=8, writedata=42, we=1 before rising edge
// (readdata should only update in asynch)
we=1;  #100;
$display("[SYNCH] Testing addr=8 with writedata=42 and we=1 (falling edge): DM[8]=2"); 
verifyEqual32(readdataSynch, 2);
///////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////
// Test: addr=8, writedata=42, we=1 after rising edge
// (Read data should update in both)
#100;
$display("[SYNCH] Testing addr=8 with writedata=42 and we=1 (falling edge): DM[8]=2"); 
verifyEqual32(readdataSynch, 42);
$display("All tests passed.");
end
///////////////////////////////////////////////////////////////////////////

endmodule